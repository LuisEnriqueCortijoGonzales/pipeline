// File pipeline_stages/execute.v

parameter ALU_FLAGS_WIDTH = 4;
parameter DATA_WIDTH = 32;

module execute (
    input wire i_clk,   // Clock signal
    input wire i_reset, // Reset signal

    input wire i_PCSource_E,
    input wire i_RegWriteEnable_E,
    input wire i_MemToReg_E,
    input wire i_MemWriteEnable_E,
    input wire [2:0] i_ALUControl_E,
    input wire i_Branch_E,
    input wire i_ALUSrc_E,
    input wire [1:0] i_FlagWrite_E,
    input wire [3:0] i_Cond_E,
    input wire [ALU_FLAGS_WIDTH-1:0] i_Flags_E,

    // Datapath
    input wire [DATA_WIDTH - 1 : 0] i_RD1_E,
    input wire [DATA_WIDTH - 1 : 0] i_RD2_E,
    input wire [DATA_WIDTH - 1 : 0] i_ExtendedImmediate_E,
    // WA3E is just pipelined

    // OUTPUTS:
    output wire [DATA_WIDTH - 1 : 0] o_Flags_E,
    output wire [DATA_WIDTH - 1 : 0] o_ALUResult_E,
    output wire [DATA_WIDTH - 1 : 0] o_WriteData_E,

    // cond unit outputs
    output reg o_PCSrc_E,
    output reg o_RegWrite_E,
    output reg o_MemToReg_E,
    output reg o_MemWrite_E
);

  wire [DATA_WIDTH - 1 : 0] SrcB_E;  // Source B for ALU
  wire ALUFlags_E[ALU_FLAGS_WIDTH - 1 : 0];  // Flags generated by ALU
  wire CondEx_E;  // Extended condition for conditional unit


  // Mux for ALU Source B: Register Data or Extended Immediate
  mux2 #(32) srcb_mux (
      .d0(i_RD2_E),
      .d1(i_EXTEndedImmediate_E),
      .s (i_ALUSrc_E),
      .y (SrcB_E)
  );

  // ALU Operations
  alu arithmetic_logic_unit (
      .a(i_RD1_E),
      .b(SrcB_E),
      .ALUControl(i_ALUControl_E),
      .Result(o_ALUResult_E),
      .ALUFlags(ALUFlags_E)
  );

  cond_unit conditional_unit (
      .i_clk(i_clk),
      .i_reset(i_reset),
      .i_FlagWrite_E(i_FlagWrite_E),
      .i_Cond_E(i_Cond_E),
      .i_Flags_E(i_Flags_E),
      .i_ALUFlags(ALUFlags_E),
      .o_Flags(o_Flags_E),
      .o_CondEx_E(CondEx_E)
  );


  wire and_1;
  wire and_2;

  assign and_1 = PCSource_E & CondEx_E;
  assign and_2 = Branch_E & CondEx_E;

  assign o_PCSrc_E = and_1 | and_2;
  assign o_RegWrite_E = i_RegWriteEnable_E & CondEx_E;
  assign o_MemToReg_E = i_MemToReg_E;
  assign o_MemWrite_E = i_MemWriteEnable_E & CondEx_E;

endmodule
