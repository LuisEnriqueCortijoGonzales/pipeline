module arm (
    input wire clk,
    input wire reset,
    output wire [31:0] PCF,
    input wire [31:0] InstrF,
    output wire MemWriteM,
    output wire [(DATA_WIDTH*2)-1:0] ALUOutM,
    output wire [31:0] WriteDataM,
    input wire [31:0] ReadDataM,
    output wire [DATA_WIDTH-1:0] R0,
    output wire [DATA_WIDTH-1:0] R1
);
  localparam ALUCONTROL_WIDTH = 6;
  localparam ALU_FLAGS_WIDTH = 5;
  parameter DATA_WIDTH = 32;

  wire [1:0] RegSrcD;
  wire [1:0] ImmSrcD;
  wire [ALUCONTROL_WIDTH-1:0] ALUControlE;
  wire ALUSrcE;
  wire BranchTakenE;
  wire MemtoRegW;
  wire [1:0] RegWriteW;
  wire [ALU_FLAGS_WIDTH-1:0] ALUFlagsE;
  wire [31:0] InstrD;
  wire [1:0] RegWriteM;
  wire MemtoRegE;
  wire PCWrPendingF;
  wire [1:0] ForwardAE;
  wire [1:0] ForwardBE;
  wire [1:0] ForwardCE;
  wire [1:0] ForwardDE;
  wire StallF;
  wire StallD;
  wire FlushD;
  wire FlushE;
  wire Match_1E_M;
  wire Match_1E_W;
  wire Match_2E_M;
  wire Match_2E_W;
  wire Match_3E_M;
  wire Match_3E_W;
  wire Match_4E_M;
  wire Match_4E_W;
  wire Match_12D_E;
  wire taken;
  //wire predict_taken;

  wire is_memory_strE;
  wire is_memory_postE;
  wire is_memory_strW;
  wire is_memory_postW;

  wire [ALU_FLAGS_WIDTH-1:0] FlagsE;
  wire [31:0] PCPlus8D;
  wire [31:0] PCPlus4F;
  wire [31:0] PredictedBranchPC;

  wire PredictTakenF;
  wire PredictTakenD;
  wire PredictTakenE;

  wire WrongPredictionE = PredictTakenE != BranchTakenE;

  wire shiftedE;

  controller Control_unit (
      .clk(clk),
      .reset(reset),
      .InstrD(InstrD[31:12]),
      .ALUFlagsE(ALUFlagsE),
      .RegSrcD(RegSrcD),
      .ImmSrcD(ImmSrcD),
      .ALUSrcE(ALUSrcE),
      .BranchTakenE(BranchTakenE),
      .PredictTakenE(PredictTakenE),
      .ALUControlE(ALUControlE),
      .MemWriteM(MemWriteM),
      .MemtoRegW(MemtoRegW),
      .RegWriteW(RegWriteW),
      .RegWriteM(RegWriteM),
      .MemtoRegE(MemtoRegE),
      .PCWrPendingF(PCWrPendingF),
      .FlushE(FlushE),
      .FlagsE(FlagsE),
      .is_memory_strE(is_memory_strE),
      .is_memory_postE(is_memory_postE),
      .is_memory_strW(is_memory_strW),
      .shiftedE(shiftedE),
      .is_memory_postW(is_memory_postW)

  );


  datapath Data_path (
      .clk(clk),
      .reset(reset),
      .RegSrcD(RegSrcD),
      .ImmSrcD(ImmSrcD),
      .ALUSrcE(ALUSrcE),
      .BranchTakenE(BranchTakenE),
      .ALUControlE(ALUControlE),
      .MemtoRegW(MemtoRegW),
      .PredictTakenF(PredictTakenF),
      .PredictedBranchPC(PredictedBranchPC),
      .RegWriteW(RegWriteW),
      .is_memory_strE(is_memory_strE),
      .is_memory_postE(is_memory_postE),
      .is_memory_strW(is_memory_strW),
      .is_memory_postW(is_memory_postW),
      .PCF(PCF),
      .InstrF(InstrF),
      .InstrD(InstrD),
      .ALUOutM(ALUOutM),
      .WriteDataM(WriteDataM),
      .ReadDataM(ReadDataM),
      .ALUFlagsE(ALUFlagsE),
      .FlagsE(FlagsE),
      .Match_1E_M(Match_1E_M),
      .Match_1E_W(Match_1E_W),
      .Match_2E_M(Match_2E_M),
      .Match_2E_W(Match_2E_W),
      .Match_3E_M(Match_3E_M),
      .Match_3E_W(Match_3E_W),
      .Match_4E_M(Match_4E_M),
      .Match_4E_W(Match_4E_W),
      .Match_12D_E(Match_12D_E),
      .ForwardAE(ForwardAE),
      .ForwardBE(ForwardBE),
      .ForwardCE(ForwardCE),
      .ForwardDE(ForwardDE),
      .StallF(StallF),
      .StallD(StallD),
      .FlushD(FlushD),
      .R0(R0),
      .R1(R1),
      .PCPlus8D(PCPlus8D),
      .PCPlus4F(PCPlus4F),
      .isBranchF(isBranchF),
      .shiftedE(shiftedE),
      .WrongPredictionE(WrongPredictionE)
  );


  // Unidad de Hazard: Detecta dependencias de datos y genera señales de control
  // para evitar conflictos en el pipeline. Maneja riesgos de datos y controla
  // el forwarding y el stalling de instrucciones.
  hazardUnit Hazard_unit (
      .clk(clk),
      .reset(reset),
      .Match_1E_M(Match_1E_M),
      .Match_1E_W(Match_1E_W),
      .Match_2E_M(Match_2E_M),
      .Match_2E_W(Match_2E_W),
      .Match_3E_M(Match_3E_M),
      .Match_3E_W(Match_3E_W),
      .Match_4E_M(Match_4E_M),
      .Match_4E_W(Match_4E_W),
      .Match_12D_E(Match_12D_E),
      .RegWriteM(RegWriteM),
      .RegWriteW(RegWriteW),
      .BranchTakenE(BranchTakenE),
      .MemtoRegE(MemtoRegE),
      .PCWrPendingF(PCWrPendingF),
      .ForwardAE(ForwardAE),
      .ForwardBE(ForwardBE),
      .ForwardCE(ForwardCE),
      .ForwardDE(ForwardDE),
      .StallF(StallF),
      .StallD(StallD),
      .FlushD(FlushD),
      .FlushE(FlushE),
      .WrongPredictionE(WrongPredictionE)
  );

  wire isBranchF = InstrF[27:26] == 2'b01;
  branch_predictor bp (
      .clk(clk),
      .reset(reset),
      .branch(isBranchF),
      .taken(BranchTakenE),
      .predict_taken(PredictTakenF)
  );
  // if ~branch, PredictTakenF = 0
  assign PredictedBranchPC = {{6{InstrF[23]}}, InstrF[23:0], 2'b00} + PCPlus4F + 4;


  // Propagate predict taken

  registro_flanco_positivo #(
      .WIDTH(1)
  ) reg_PredictTaken_FD (
      .clk(clk),  // Reloj del sistema
      .reset(reset),  // Señal de reinicio
      .d(PredictTakenF),  // Dato de entrada
      .q(PredictTakenD)  // Dato de salida
  );


  registro_flanco_positivo_habilitacion_limpieza #(
      .WIDTH(1)
  ) reg_PredictTaken_DE (
      .clk(clk),
      .reset(reset),
      .en(1'b1),
      .clear(FlushE),
      .clear_value(1'b0),
      .d(PredictTakenD),
      .q(PredictTakenE)
  );


endmodule
