// File: datapath.v
module datapath (
    clk,
    reset
);

  input clk;
  input reset;


  // FETCH


endmodule
